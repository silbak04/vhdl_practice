--===========================================================================--
--===============================  VHDL  ====================================--
--===========================================================================--
--                                                                           --
-- FILE NAME:     full_adder.vhd                                             --
--                                                                           --
-- DATE:          4/12/2011                                                  --
--                                                                           --
-- DESIGNER:      Samir Silbak                                               --
--                                                                           --
-- DESCRIPTION:   1-bit full adder                                           --
--                                                                           --
--===========================================================================--
--===============================  VHDL  ====================================--
--===========================================================================--

library ieee;
library work;
use ieee.std_logic_1164.all;

--===========================================================================--
--===============================  I/O Ports  ===============================--
--===========================================================================--

entity full_adder is
    port(
        a           : in  std_logic;
        b           : in  std_logic;
        cin         : in  std_logic;
        s           : out std_logic;
        cout        : out std_logic
    );
end full_adder;

--===========================================================================--
--=============================  Main Function  =============================--
--===========================================================================--

architecture data_flow of full_adder is
begin

    s <= a xor b xor cin;
    cout <= (a and b) or (a and cin) or
            (b and cin);

end data_flow;
